VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_wishbone_demo
  CLASS BLOCK ;
  FOREIGN wrapped_wishbone_demo ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 220.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 95.240 100.000 95.840 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 68.040 100.000 68.640 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 61.240 100.000 61.840 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 131.960 100.000 132.560 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 107.480 100.000 108.080 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 4.120 100.000 4.720 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 216.000 13.250 220.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 44.920 100.000 45.520 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 171.400 100.000 172.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 216.000 81.330 220.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 216.000 89.610 220.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 216.000 33.490 220.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 216.000 6.810 220.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 47.640 100.000 48.240 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 100.680 100.000 101.280 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 161.880 100.000 162.480 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 10.920 100.000 11.520 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 8.200 100.000 8.800 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 216.000 64.770 220.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 17.720 100.000 18.320 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 216.000 69.370 220.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 148.280 100.000 148.880 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 185.000 100.000 185.600 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 144.200 100.000 144.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 216.000 87.770 220.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 51.720 100.000 52.320 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 204.040 100.000 204.640 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 216.000 76.730 220.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 141.480 100.000 142.080 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 216.000 31.650 220.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 216.000 96.970 220.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 216.000 44.530 220.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 194.520 100.000 195.120 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 198.600 100.000 199.200 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 216.000 78.570 220.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 155.080 100.000 155.680 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 91.160 100.000 91.760 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 208.120 100.000 208.720 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 127.880 100.000 128.480 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 216.000 51.890 220.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 216.000 98.810 220.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 216.000 19.690 220.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 81.640 100.000 82.240 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 216.000 83.170 220.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 15.000 100.000 15.600 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 216.000 94.210 220.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 216.000 58.330 220.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 151.000 100.000 151.600 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 38.120 100.000 38.720 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 118.360 100.000 118.960 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 216.000 49.130 220.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 216.000 67.530 220.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 97.960 100.000 98.560 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 216.000 56.490 220.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 216.000 4.050 220.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 216.000 24.290 220.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 216.000 42.690 220.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 34.040 100.000 34.640 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 54.440 100.000 55.040 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 216.000 40.850 220.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 121.080 100.000 121.680 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 74.840 100.000 75.440 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 191.800 100.000 192.400 ;
    END
  END io_out[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.545 10.640 21.145 206.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.195 10.640 50.795 206.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.850 10.640 80.450 206.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 34.370 10.640 35.970 206.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.025 10.640 65.625 206.960 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 216.000 16.010 220.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 214.920 100.000 215.520 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 157.800 100.000 158.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 187.720 100.000 188.320 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 84.360 100.000 84.960 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 216.000 38.090 220.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 70.760 100.000 71.360 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 31.320 100.000 31.920 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 137.400 100.000 138.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 24.520 100.000 25.120 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 216.000 11.410 220.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 216.000 8.650 220.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 58.520 100.000 59.120 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 180.920 100.000 181.520 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 1.400 100.000 2.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 216.000 73.970 220.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 216.000 2.210 220.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 216.000 22.450 220.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 216.000 17.850 220.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 210.840 100.000 211.440 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 216.000 36.250 220.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 104.760 100.000 105.360 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 174.120 100.000 174.720 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 134.680 100.000 135.280 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 201.320 100.000 201.920 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 216.000 47.290 220.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 111.560 100.000 112.160 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 63.960 100.000 64.560 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 21.800 100.000 22.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 88.440 100.000 89.040 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 217.640 100.000 218.240 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 27.240 100.000 27.840 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 114.280 100.000 114.880 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 178.200 100.000 178.800 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 216.000 92.370 220.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 40.840 100.000 41.440 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 216.000 85.930 220.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 216.000 28.890 220.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 216.000 53.730 220.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 216.000 27.050 220.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 216.000 72.130 220.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 77.560 100.000 78.160 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 167.320 100.000 167.920 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 164.600 100.000 165.200 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 216.000 62.930 220.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 216.000 61.090 220.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 125.160 100.000 125.760 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 95.535 215.135 ;
      LAYER met1 ;
        RECT 0.070 10.640 98.830 215.180 ;
      LAYER met2 ;
        RECT 0.100 215.720 1.650 219.485 ;
        RECT 2.490 215.720 3.490 219.485 ;
        RECT 4.330 215.720 6.250 219.485 ;
        RECT 7.090 215.720 8.090 219.485 ;
        RECT 8.930 215.720 10.850 219.485 ;
        RECT 11.690 215.720 12.690 219.485 ;
        RECT 13.530 215.720 15.450 219.485 ;
        RECT 16.290 215.720 17.290 219.485 ;
        RECT 18.130 215.720 19.130 219.485 ;
        RECT 19.970 215.720 21.890 219.485 ;
        RECT 22.730 215.720 23.730 219.485 ;
        RECT 24.570 215.720 26.490 219.485 ;
        RECT 27.330 215.720 28.330 219.485 ;
        RECT 29.170 215.720 31.090 219.485 ;
        RECT 31.930 215.720 32.930 219.485 ;
        RECT 33.770 215.720 35.690 219.485 ;
        RECT 36.530 215.720 37.530 219.485 ;
        RECT 38.370 215.720 40.290 219.485 ;
        RECT 41.130 215.720 42.130 219.485 ;
        RECT 42.970 215.720 43.970 219.485 ;
        RECT 44.810 215.720 46.730 219.485 ;
        RECT 47.570 215.720 48.570 219.485 ;
        RECT 49.410 215.720 51.330 219.485 ;
        RECT 52.170 215.720 53.170 219.485 ;
        RECT 54.010 215.720 55.930 219.485 ;
        RECT 56.770 215.720 57.770 219.485 ;
        RECT 58.610 215.720 60.530 219.485 ;
        RECT 61.370 215.720 62.370 219.485 ;
        RECT 63.210 215.720 64.210 219.485 ;
        RECT 65.050 215.720 66.970 219.485 ;
        RECT 67.810 215.720 68.810 219.485 ;
        RECT 69.650 215.720 71.570 219.485 ;
        RECT 72.410 215.720 73.410 219.485 ;
        RECT 74.250 215.720 76.170 219.485 ;
        RECT 77.010 215.720 78.010 219.485 ;
        RECT 78.850 215.720 80.770 219.485 ;
        RECT 81.610 215.720 82.610 219.485 ;
        RECT 83.450 215.720 85.370 219.485 ;
        RECT 86.210 215.720 87.210 219.485 ;
        RECT 88.050 215.720 89.050 219.485 ;
        RECT 89.890 215.720 91.810 219.485 ;
        RECT 92.650 215.720 93.650 219.485 ;
        RECT 94.490 215.720 96.410 219.485 ;
        RECT 97.250 215.720 98.250 219.485 ;
        RECT 0.100 4.280 98.800 215.720 ;
        RECT 0.650 1.515 1.650 4.280 ;
        RECT 2.490 1.515 3.490 4.280 ;
        RECT 4.330 1.515 6.250 4.280 ;
        RECT 7.090 1.515 8.090 4.280 ;
        RECT 8.930 1.515 10.850 4.280 ;
        RECT 11.690 1.515 12.690 4.280 ;
        RECT 13.530 1.515 15.450 4.280 ;
        RECT 16.290 1.515 17.290 4.280 ;
        RECT 18.130 1.515 20.050 4.280 ;
        RECT 20.890 1.515 21.890 4.280 ;
        RECT 22.730 1.515 23.730 4.280 ;
        RECT 24.570 1.515 26.490 4.280 ;
        RECT 27.330 1.515 28.330 4.280 ;
        RECT 29.170 1.515 31.090 4.280 ;
        RECT 31.930 1.515 32.930 4.280 ;
        RECT 33.770 1.515 35.690 4.280 ;
        RECT 36.530 1.515 37.530 4.280 ;
        RECT 38.370 1.515 40.290 4.280 ;
        RECT 41.130 1.515 42.130 4.280 ;
        RECT 42.970 1.515 44.890 4.280 ;
        RECT 45.730 1.515 46.730 4.280 ;
        RECT 47.570 1.515 48.570 4.280 ;
        RECT 49.410 1.515 51.330 4.280 ;
        RECT 52.170 1.515 53.170 4.280 ;
        RECT 54.010 1.515 55.930 4.280 ;
        RECT 56.770 1.515 57.770 4.280 ;
        RECT 58.610 1.515 60.530 4.280 ;
        RECT 61.370 1.515 62.370 4.280 ;
        RECT 63.210 1.515 65.130 4.280 ;
        RECT 65.970 1.515 66.970 4.280 ;
        RECT 67.810 1.515 69.730 4.280 ;
        RECT 70.570 1.515 71.570 4.280 ;
        RECT 72.410 1.515 73.410 4.280 ;
        RECT 74.250 1.515 76.170 4.280 ;
        RECT 77.010 1.515 78.010 4.280 ;
        RECT 78.850 1.515 80.770 4.280 ;
        RECT 81.610 1.515 82.610 4.280 ;
        RECT 83.450 1.515 85.370 4.280 ;
        RECT 86.210 1.515 87.210 4.280 ;
        RECT 88.050 1.515 89.970 4.280 ;
        RECT 90.810 1.515 91.810 4.280 ;
        RECT 92.650 1.515 94.570 4.280 ;
        RECT 95.410 1.515 96.410 4.280 ;
        RECT 97.250 1.515 98.250 4.280 ;
      LAYER met3 ;
        RECT 4.400 218.640 96.000 219.465 ;
        RECT 4.400 218.600 95.600 218.640 ;
        RECT 4.000 217.280 95.600 218.600 ;
        RECT 4.400 217.240 95.600 217.280 ;
        RECT 4.400 215.920 96.000 217.240 ;
        RECT 4.400 215.880 95.600 215.920 ;
        RECT 4.000 214.520 95.600 215.880 ;
        RECT 4.000 213.200 96.000 214.520 ;
        RECT 4.400 211.840 96.000 213.200 ;
        RECT 4.400 211.800 95.600 211.840 ;
        RECT 4.000 210.480 95.600 211.800 ;
        RECT 4.400 210.440 95.600 210.480 ;
        RECT 4.400 209.120 96.000 210.440 ;
        RECT 4.400 209.080 95.600 209.120 ;
        RECT 4.000 207.760 95.600 209.080 ;
        RECT 4.400 207.720 95.600 207.760 ;
        RECT 4.400 206.360 96.000 207.720 ;
        RECT 4.000 205.040 96.000 206.360 ;
        RECT 4.000 203.680 95.600 205.040 ;
        RECT 4.400 203.640 95.600 203.680 ;
        RECT 4.400 202.320 96.000 203.640 ;
        RECT 4.400 202.280 95.600 202.320 ;
        RECT 4.000 200.960 95.600 202.280 ;
        RECT 4.400 200.920 95.600 200.960 ;
        RECT 4.400 199.600 96.000 200.920 ;
        RECT 4.400 199.560 95.600 199.600 ;
        RECT 4.000 198.200 95.600 199.560 ;
        RECT 4.000 196.880 96.000 198.200 ;
        RECT 4.400 195.520 96.000 196.880 ;
        RECT 4.400 195.480 95.600 195.520 ;
        RECT 4.000 194.160 95.600 195.480 ;
        RECT 4.400 194.120 95.600 194.160 ;
        RECT 4.400 192.800 96.000 194.120 ;
        RECT 4.400 192.760 95.600 192.800 ;
        RECT 4.000 191.400 95.600 192.760 ;
        RECT 4.000 190.080 96.000 191.400 ;
        RECT 4.400 188.720 96.000 190.080 ;
        RECT 4.400 188.680 95.600 188.720 ;
        RECT 4.000 187.360 95.600 188.680 ;
        RECT 4.400 187.320 95.600 187.360 ;
        RECT 4.400 186.000 96.000 187.320 ;
        RECT 4.400 185.960 95.600 186.000 ;
        RECT 4.000 184.600 95.600 185.960 ;
        RECT 4.000 183.280 96.000 184.600 ;
        RECT 4.400 181.920 96.000 183.280 ;
        RECT 4.400 181.880 95.600 181.920 ;
        RECT 4.000 180.560 95.600 181.880 ;
        RECT 4.400 180.520 95.600 180.560 ;
        RECT 4.400 179.200 96.000 180.520 ;
        RECT 4.400 179.160 95.600 179.200 ;
        RECT 4.000 177.800 95.600 179.160 ;
        RECT 4.000 176.480 96.000 177.800 ;
        RECT 4.400 175.120 96.000 176.480 ;
        RECT 4.400 175.080 95.600 175.120 ;
        RECT 4.000 173.760 95.600 175.080 ;
        RECT 4.400 173.720 95.600 173.760 ;
        RECT 4.400 172.400 96.000 173.720 ;
        RECT 4.400 172.360 95.600 172.400 ;
        RECT 4.000 171.040 95.600 172.360 ;
        RECT 4.400 171.000 95.600 171.040 ;
        RECT 4.400 169.640 96.000 171.000 ;
        RECT 4.000 168.320 96.000 169.640 ;
        RECT 4.000 166.960 95.600 168.320 ;
        RECT 4.400 166.920 95.600 166.960 ;
        RECT 4.400 165.600 96.000 166.920 ;
        RECT 4.400 165.560 95.600 165.600 ;
        RECT 4.000 164.240 95.600 165.560 ;
        RECT 4.400 164.200 95.600 164.240 ;
        RECT 4.400 162.880 96.000 164.200 ;
        RECT 4.400 162.840 95.600 162.880 ;
        RECT 4.000 161.480 95.600 162.840 ;
        RECT 4.000 160.160 96.000 161.480 ;
        RECT 4.400 158.800 96.000 160.160 ;
        RECT 4.400 158.760 95.600 158.800 ;
        RECT 4.000 157.440 95.600 158.760 ;
        RECT 4.400 157.400 95.600 157.440 ;
        RECT 4.400 156.080 96.000 157.400 ;
        RECT 4.400 156.040 95.600 156.080 ;
        RECT 4.000 154.680 95.600 156.040 ;
        RECT 4.000 153.360 96.000 154.680 ;
        RECT 4.400 152.000 96.000 153.360 ;
        RECT 4.400 151.960 95.600 152.000 ;
        RECT 4.000 150.640 95.600 151.960 ;
        RECT 4.400 150.600 95.600 150.640 ;
        RECT 4.400 149.280 96.000 150.600 ;
        RECT 4.400 149.240 95.600 149.280 ;
        RECT 4.000 147.880 95.600 149.240 ;
        RECT 4.000 146.560 96.000 147.880 ;
        RECT 4.400 145.200 96.000 146.560 ;
        RECT 4.400 145.160 95.600 145.200 ;
        RECT 4.000 143.840 95.600 145.160 ;
        RECT 4.400 143.800 95.600 143.840 ;
        RECT 4.400 142.480 96.000 143.800 ;
        RECT 4.400 142.440 95.600 142.480 ;
        RECT 4.000 141.120 95.600 142.440 ;
        RECT 4.400 141.080 95.600 141.120 ;
        RECT 4.400 139.720 96.000 141.080 ;
        RECT 4.000 138.400 96.000 139.720 ;
        RECT 4.000 137.040 95.600 138.400 ;
        RECT 4.400 137.000 95.600 137.040 ;
        RECT 4.400 135.680 96.000 137.000 ;
        RECT 4.400 135.640 95.600 135.680 ;
        RECT 4.000 134.320 95.600 135.640 ;
        RECT 4.400 134.280 95.600 134.320 ;
        RECT 4.400 132.960 96.000 134.280 ;
        RECT 4.400 132.920 95.600 132.960 ;
        RECT 4.000 131.560 95.600 132.920 ;
        RECT 4.000 130.240 96.000 131.560 ;
        RECT 4.400 128.880 96.000 130.240 ;
        RECT 4.400 128.840 95.600 128.880 ;
        RECT 4.000 127.520 95.600 128.840 ;
        RECT 4.400 127.480 95.600 127.520 ;
        RECT 4.400 126.160 96.000 127.480 ;
        RECT 4.400 126.120 95.600 126.160 ;
        RECT 4.000 124.760 95.600 126.120 ;
        RECT 4.000 123.440 96.000 124.760 ;
        RECT 4.400 122.080 96.000 123.440 ;
        RECT 4.400 122.040 95.600 122.080 ;
        RECT 4.000 120.720 95.600 122.040 ;
        RECT 4.400 120.680 95.600 120.720 ;
        RECT 4.400 119.360 96.000 120.680 ;
        RECT 4.400 119.320 95.600 119.360 ;
        RECT 4.000 117.960 95.600 119.320 ;
        RECT 4.000 116.640 96.000 117.960 ;
        RECT 4.400 115.280 96.000 116.640 ;
        RECT 4.400 115.240 95.600 115.280 ;
        RECT 4.000 113.920 95.600 115.240 ;
        RECT 4.400 113.880 95.600 113.920 ;
        RECT 4.400 112.560 96.000 113.880 ;
        RECT 4.400 112.520 95.600 112.560 ;
        RECT 4.000 111.160 95.600 112.520 ;
        RECT 4.000 109.840 96.000 111.160 ;
        RECT 4.400 108.480 96.000 109.840 ;
        RECT 4.400 108.440 95.600 108.480 ;
        RECT 4.000 107.120 95.600 108.440 ;
        RECT 4.400 107.080 95.600 107.120 ;
        RECT 4.400 105.760 96.000 107.080 ;
        RECT 4.400 105.720 95.600 105.760 ;
        RECT 4.000 104.400 95.600 105.720 ;
        RECT 4.400 104.360 95.600 104.400 ;
        RECT 4.400 103.000 96.000 104.360 ;
        RECT 4.000 101.680 96.000 103.000 ;
        RECT 4.000 100.320 95.600 101.680 ;
        RECT 4.400 100.280 95.600 100.320 ;
        RECT 4.400 98.960 96.000 100.280 ;
        RECT 4.400 98.920 95.600 98.960 ;
        RECT 4.000 97.600 95.600 98.920 ;
        RECT 4.400 97.560 95.600 97.600 ;
        RECT 4.400 96.240 96.000 97.560 ;
        RECT 4.400 96.200 95.600 96.240 ;
        RECT 4.000 94.840 95.600 96.200 ;
        RECT 4.000 93.520 96.000 94.840 ;
        RECT 4.400 92.160 96.000 93.520 ;
        RECT 4.400 92.120 95.600 92.160 ;
        RECT 4.000 90.800 95.600 92.120 ;
        RECT 4.400 90.760 95.600 90.800 ;
        RECT 4.400 89.440 96.000 90.760 ;
        RECT 4.400 89.400 95.600 89.440 ;
        RECT 4.000 88.040 95.600 89.400 ;
        RECT 4.000 86.720 96.000 88.040 ;
        RECT 4.400 85.360 96.000 86.720 ;
        RECT 4.400 85.320 95.600 85.360 ;
        RECT 4.000 84.000 95.600 85.320 ;
        RECT 4.400 83.960 95.600 84.000 ;
        RECT 4.400 82.640 96.000 83.960 ;
        RECT 4.400 82.600 95.600 82.640 ;
        RECT 4.000 81.240 95.600 82.600 ;
        RECT 4.000 79.920 96.000 81.240 ;
        RECT 4.400 78.560 96.000 79.920 ;
        RECT 4.400 78.520 95.600 78.560 ;
        RECT 4.000 77.200 95.600 78.520 ;
        RECT 4.400 77.160 95.600 77.200 ;
        RECT 4.400 75.840 96.000 77.160 ;
        RECT 4.400 75.800 95.600 75.840 ;
        RECT 4.000 74.440 95.600 75.800 ;
        RECT 4.000 73.120 96.000 74.440 ;
        RECT 4.400 71.760 96.000 73.120 ;
        RECT 4.400 71.720 95.600 71.760 ;
        RECT 4.000 70.400 95.600 71.720 ;
        RECT 4.400 70.360 95.600 70.400 ;
        RECT 4.400 69.040 96.000 70.360 ;
        RECT 4.400 69.000 95.600 69.040 ;
        RECT 4.000 67.680 95.600 69.000 ;
        RECT 4.400 67.640 95.600 67.680 ;
        RECT 4.400 66.280 96.000 67.640 ;
        RECT 4.000 64.960 96.000 66.280 ;
        RECT 4.000 63.600 95.600 64.960 ;
        RECT 4.400 63.560 95.600 63.600 ;
        RECT 4.400 62.240 96.000 63.560 ;
        RECT 4.400 62.200 95.600 62.240 ;
        RECT 4.000 60.880 95.600 62.200 ;
        RECT 4.400 60.840 95.600 60.880 ;
        RECT 4.400 59.520 96.000 60.840 ;
        RECT 4.400 59.480 95.600 59.520 ;
        RECT 4.000 58.120 95.600 59.480 ;
        RECT 4.000 56.800 96.000 58.120 ;
        RECT 4.400 55.440 96.000 56.800 ;
        RECT 4.400 55.400 95.600 55.440 ;
        RECT 4.000 54.080 95.600 55.400 ;
        RECT 4.400 54.040 95.600 54.080 ;
        RECT 4.400 52.720 96.000 54.040 ;
        RECT 4.400 52.680 95.600 52.720 ;
        RECT 4.000 51.320 95.600 52.680 ;
        RECT 4.000 50.000 96.000 51.320 ;
        RECT 4.400 48.640 96.000 50.000 ;
        RECT 4.400 48.600 95.600 48.640 ;
        RECT 4.000 47.280 95.600 48.600 ;
        RECT 4.400 47.240 95.600 47.280 ;
        RECT 4.400 45.920 96.000 47.240 ;
        RECT 4.400 45.880 95.600 45.920 ;
        RECT 4.000 44.520 95.600 45.880 ;
        RECT 4.000 43.200 96.000 44.520 ;
        RECT 4.400 41.840 96.000 43.200 ;
        RECT 4.400 41.800 95.600 41.840 ;
        RECT 4.000 40.480 95.600 41.800 ;
        RECT 4.400 40.440 95.600 40.480 ;
        RECT 4.400 39.120 96.000 40.440 ;
        RECT 4.400 39.080 95.600 39.120 ;
        RECT 4.000 37.720 95.600 39.080 ;
        RECT 4.000 36.400 96.000 37.720 ;
        RECT 4.400 35.040 96.000 36.400 ;
        RECT 4.400 35.000 95.600 35.040 ;
        RECT 4.000 33.680 95.600 35.000 ;
        RECT 4.400 33.640 95.600 33.680 ;
        RECT 4.400 32.320 96.000 33.640 ;
        RECT 4.400 32.280 95.600 32.320 ;
        RECT 4.000 30.960 95.600 32.280 ;
        RECT 4.400 30.920 95.600 30.960 ;
        RECT 4.400 29.560 96.000 30.920 ;
        RECT 4.000 28.240 96.000 29.560 ;
        RECT 4.000 26.880 95.600 28.240 ;
        RECT 4.400 26.840 95.600 26.880 ;
        RECT 4.400 25.520 96.000 26.840 ;
        RECT 4.400 25.480 95.600 25.520 ;
        RECT 4.000 24.160 95.600 25.480 ;
        RECT 4.400 24.120 95.600 24.160 ;
        RECT 4.400 22.800 96.000 24.120 ;
        RECT 4.400 22.760 95.600 22.800 ;
        RECT 4.000 21.400 95.600 22.760 ;
        RECT 4.000 20.080 96.000 21.400 ;
        RECT 4.400 18.720 96.000 20.080 ;
        RECT 4.400 18.680 95.600 18.720 ;
        RECT 4.000 17.360 95.600 18.680 ;
        RECT 4.400 17.320 95.600 17.360 ;
        RECT 4.400 16.000 96.000 17.320 ;
        RECT 4.400 15.960 95.600 16.000 ;
        RECT 4.000 14.600 95.600 15.960 ;
        RECT 4.000 13.280 96.000 14.600 ;
        RECT 4.400 11.920 96.000 13.280 ;
        RECT 4.400 11.880 95.600 11.920 ;
        RECT 4.000 10.560 95.600 11.880 ;
        RECT 4.400 10.520 95.600 10.560 ;
        RECT 4.400 9.200 96.000 10.520 ;
        RECT 4.400 9.160 95.600 9.200 ;
        RECT 4.000 7.800 95.600 9.160 ;
        RECT 4.000 6.480 96.000 7.800 ;
        RECT 4.400 5.120 96.000 6.480 ;
        RECT 4.400 5.080 95.600 5.120 ;
        RECT 4.000 3.760 95.600 5.080 ;
        RECT 4.400 3.720 95.600 3.760 ;
        RECT 4.400 2.400 96.000 3.720 ;
        RECT 4.400 2.360 95.600 2.400 ;
        RECT 4.000 1.535 95.600 2.360 ;
      LAYER met4 ;
        RECT 51.195 10.640 52.145 206.960 ;
  END
END wrapped_wishbone_demo
END LIBRARY

